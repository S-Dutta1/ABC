// Benchmark "file" written by ABC on Tue Nov 29 19:02:41 2016

module file ( 
    a, b, c, d,
    f3  );
  input  a, b, c, d;
  output f3;
  assign f3 = a ^ ~b;
endmodule


